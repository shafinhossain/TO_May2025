* Extracted by KLayout with SG13G2 LVS runset on : 12/05/2025 06:49

.SUBCKT FMD_QNC_10_8way_PA_180G RFIN|RFOUT|VSS VCC1 VBB2 VCC2 VBB1 VCC2$1 VCC1$1
Q$1 \$82446 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$21 \$83131 \$85521 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$39 \$84298 \$85326 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$57 \$131269 \$133283 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$75 \$132284 \$134518 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$93 \$133085 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$113 \$221730 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$133 \$222590 \$225693 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$151 \$223429 \$226742 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$169 \$271505 \$273222 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$187 \$272424 \$273416 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$205 \$272822 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$225 \$364675 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$245 \$365713 \$366748 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$263 \$366747 \$367591 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$281 \$414487 \$416346 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$299 \$415359 \$417246 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$317 \$415756 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$337 \$505016 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$357 \$505608 \$508035 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$375 \$506607 \$507841 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$393 \$554728 \$555602 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$411 \$555603 \$557289 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=57.1475p PB=41.52u AC=57.123234p PC=41.51u NE=18 m=18
Q$429 \$556037 RFIN|RFOUT|VSS RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
R$449 RFIN|RFOUT|VSS VBB2 rsil w=2u l=12u ps=0 b=0 m=8
R$450 \$85521 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$451 \$85326 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$452 RFIN|RFOUT|VSS RFIN|RFOUT|VSS rsil w=2.04u l=28u ps=0 b=0 m=14
R$454 VBB1 \$133283 rsil w=2u l=11u ps=0 b=0 m=1
R$455 VBB1 \$134518 rsil w=2u l=11u ps=0 b=0 m=1
R$460 \$225693 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$461 \$226742 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$464 VBB1 \$273222 rsil w=2u l=11u ps=0 b=0 m=1
R$465 VBB1 \$273416 rsil w=2u l=11u ps=0 b=0 m=1
R$470 \$366748 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$471 \$367591 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$474 VBB1 \$416346 rsil w=2u l=11u ps=0 b=0 m=1
R$475 VBB1 \$417246 rsil w=2u l=11u ps=0 b=0 m=1
R$480 \$508035 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$481 \$507841 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$484 VBB1 \$555602 rsil w=2u l=11u ps=0 b=0 m=1
R$485 VBB1 \$557289 rsil w=2u l=11u ps=0 b=0 m=1
R$487 VCC2 \$82446 rppd w=35u l=2u ps=0 b=0 m=1
R$488 VCC1 \$83131 rppd w=35u l=2u ps=0 b=0 m=1
R$489 VCC1 \$84298 rppd w=35u l=2u ps=0 b=0 m=1
R$490 \$131269 VCC1 rppd w=35u l=2u ps=0 b=0 m=1
R$491 \$132284 VCC1 rppd w=35u l=2u ps=0 b=0 m=1
R$492 \$133085 VCC2 rppd w=35u l=2u ps=0 b=0 m=1
R$493 VCC2 \$221730 rppd w=35u l=2u ps=0 b=0 m=1
R$494 VCC1 \$222590 rppd w=35u l=2u ps=0 b=0 m=1
R$495 VCC1 \$223429 rppd w=35u l=2u ps=0 b=0 m=1
R$496 \$271505 VCC1 rppd w=35u l=2u ps=0 b=0 m=1
R$497 \$272424 VCC1 rppd w=35u l=2u ps=0 b=0 m=1
R$498 \$272822 VCC2$1 rppd w=35u l=2u ps=0 b=0 m=1
R$499 VCC2$1 \$364675 rppd w=35u l=2u ps=0 b=0 m=1
R$500 VCC1 \$365713 rppd w=35u l=2u ps=0 b=0 m=1
R$501 VCC1 \$366747 rppd w=35u l=2u ps=0 b=0 m=1
R$502 \$414487 VCC1$1 rppd w=35u l=2u ps=0 b=0 m=1
R$503 \$415359 VCC1$1 rppd w=35u l=2u ps=0 b=0 m=1
R$504 \$415756 VCC2$1 rppd w=35u l=2u ps=0 b=0 m=1
R$505 VCC2$1 \$505016 rppd w=35u l=2u ps=0 b=0 m=1
R$506 VCC1$1 \$505608 rppd w=35u l=2u ps=0 b=0 m=1
R$507 VCC1$1 \$506607 rppd w=35u l=2u ps=0 b=0 m=1
R$508 \$554728 VCC1$1 rppd w=35u l=2u ps=0 b=0 m=1
R$509 \$555603 VCC1$1 rppd w=35u l=2u ps=0 b=0 m=1
R$510 \$556037 VCC2$1 rppd w=35u l=2u ps=0 b=0 m=1
C$511 VCC2 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=10
C$513 VCC1 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=28
C$547 VCC2$1 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=16
C$555 VCC1$1 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=16
.ENDS FMD_QNC_10_8way_PA_180G
